module BCD2SEG (P, X, SSD);
       input [3:0] X;
		 input P;
       output [0:6] SSD;
       assign SSD[0] = (((~X[3] & ~X[2] & ~X[1] &  X[0]) | (~X[3] &  X[2] & ~X[1] & ~X[0]))) & P;
       assign SSD[1] = (((~X[3] &  X[2] & ~X[1] &  X[0]) | (~X[3] &  X[2] &  X[1] & ~X[0]))) & P;
       assign SSD[2] =  ((~X[3] & ~X[2] &  X[1] & ~X[0])) & P;
       assign SSD[3] = (((~X[3] & ~X[2] & ~X[1] &  X[0]) | (~X[3] &  X[2] & ~X[1] & ~X[0]) | (~X[3] &  X[2] & X[1] & X[0]) | (X[3] & ~X[2] & ~X[1] & X[0]))) & P;
       assign SSD[4] = (~((~X[2] & ~X[0]) | (X[1] & ~X[0]))) & P;
       assign SSD[5] = (((~X[3] & ~X[2] & ~X[1] &  X[0]) | (~X[3] & ~X[2] &  X[1] & ~X[0]) | (~X[3] & ~X[2] & X[1] & X[0]) | (~X[3] & X[2] & X[1] & X[0]))) & P;
       assign SSD[6] = (((~X[3] & ~X[2] & ~X[1] &  X[0]) | (~X[3] & ~X[2] & ~X[1] & ~X[0]) | (~X[3] &  X[2] & X[1] & X[0]))) & P;
endmodule